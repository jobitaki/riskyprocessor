parameter logic ADDR_WIDTH = 9;
parameter logic SIM_MEM_SIZE = 16'hFFFF;

typedef enum logic [4:0] {
  LB  = 32'b????????????_?????_000_?????_0000011,
  ADD = 32'b0000000_?????_?????_000_?????_0110011
} opcode_t;
