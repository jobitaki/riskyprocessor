`default_nettype none

module alu (
    input  logic [31:0] alu_in_1,
    input  logic [31:0] alu_in_2,
    input  logic [ 4:0] alu_op_sel,
    output logic [31:0] alu_out
);



endmodule : alu
