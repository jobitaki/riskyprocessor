`default_nettype none

module risky();

  // ALU + MUXES
  // REGFILE
  // MDR, MAR
  // DECODER
  // IR
  // PC

endmodule : risky
