parameter int ADDR_WIDTH = 9;
parameter int SIM_MEM_SIZE = 16'hFFFF;

typedef enum logic [31:0] {
  LB  = 32'b????_????_????_????_?000_????_?000_0011,
  ADD = 32'b0000_000?_????_????_?000_????_?011_0011
} opcode_e;
