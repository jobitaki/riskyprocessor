`default_nettype none

module execute (
  input logic [31:0] instr
);


  
endmodule : execute