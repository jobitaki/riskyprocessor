parameter int ADDR_WIDTH = 9;
parameter int SIM_MEM_SIZE = 16'hFFFF;

typedef enum logic [31:0] {
  // I-type instructions
  I_LB          = 32'b????_????_????_????_?000_????_?000_0011,
  I_LH          = 32'b????_????_????_????_?001_????_?000_0011,
  I_LW          = 32'b????_????_????_????_?010_????_?000_0011,
  I_LBU         = 32'b????_????_????_????_?100_????_?000_0011,
  I_LHU         = 32'b????_????_????_????_?101_????_?000_0011,
  I_ALL_LOADS   = 32'b????_????_????_????_????_????_?000_0011,

  // R-type instructions
  R_ADD_SUB = 32'b0?00_000?_????_????_?000_????_?011_0011,
  R_SLL     = 32'b0000_000?_????_????_?001_????_?011_0011,
  R_SLT     = 32'b0000_000?_????_????_?010_????_?011_0011,
  R_SLTU    = 32'b0000_000?_????_????_?011_????_?011_0011,
  R_XOR     = 32'b0000_000?_????_????_?100_????_?011_0011,
  R_ALL     = 32'b????_????_????_????_????_????_?011_0011
} opcode_e;

typedef enum logic [4:0] {
  ALU_ADD   = 5'b00000,
  ALU_SLL   = 5'b00001,
  ALU_SLT   = 5'b00010,
  ALU_SLTU  = 5'b00011,
  ALU_XOR   = 5'b00100,
  ALU_UNDEF = 5'b11111
} alu_op_e;
