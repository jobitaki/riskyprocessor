parameter int ADDR_WIDTH = 9;
parameter int SIM_MEM_SIZE = 16'hFFFF;

typedef enum logic [31:0] {
  // I-type instructions
  I_LB        = 32'b????_????_????_????_?000_????_?000_0011,
  I_LH        = 32'b????_????_????_????_?001_????_?000_0011,
  I_LW        = 32'b????_????_????_????_?010_????_?000_0011,
  I_LBU       = 32'b????_????_????_????_?100_????_?000_0011,
  I_LHU       = 32'b????_????_????_????_?101_????_?000_0011,
  I_ALL_LOADS = 32'b????_????_????_????_????_????_?000_0011,

  // R-type instructions
  R_ADD     = 32'b0000_000?_????_????_?000_????_?011_0011,
  R_SUB     = 32'b0100_000?_????_????_?000_????_?011_0011,
  R_SLL     = 32'b0000_000?_????_????_?001_????_?011_0011,
  R_SLT     = 32'b0000_000?_????_????_?010_????_?011_0011,
  R_SLTU    = 32'b0000_000?_????_????_?011_????_?011_0011,
  R_XOR     = 32'b0000_000?_????_????_?100_????_?011_0011,
  R_SRL     = 32'b0000_000?_????_????_?101_????_?011_0011,
  R_SRA     = 32'b0100_000?_????_????_?101_????_?011_0011,
  R_OR      = 32'b0000_000?_????_????_?110_????_?011_0011,
  R_AND     = 32'b0000_000?_????_????_?111_????_?011_0011,
  R_ALL     = 32'b????_????_????_????_????_????_?011_0011,

  // S-type instructions
  S_SB  = 32'b????_????_????_????_?000_????_?010_0011, 
  S_SH  = 32'b????_????_????_????_?001_????_?010_0011, 
  S_SW  = 32'b????_????_????_????_?010_????_?010_0011,
  S_ALL = 32'b????_????_????_????_????_????_?010_0011,

  // B-type instructions
  B_BEQ,
  B_BNE,
  B_BGE,
  B_BLTU,
  B_BGEU
} opcode_e;

typedef enum logic [4:0] {
  ALU_ADD   = 5'b00000,
  ALU_SUB   = 5'b00001,
  ALU_SLL   = 5'b00010,
  ALU_SLT   = 5'b00011,
  ALU_SLTU  = 5'b00100,
  ALU_XOR   = 5'b00101,
  ALU_SRL   = 5'b00110,
  ALU_SRA   = 5'b00111,
  ALU_OR    = 5'b01000,
  ALU_AND   = 5'b01001,
  ALU_UNDEF = 5'b11111
} alu_op_e;

typedef enum logic [1:0] {
  FU_SRC_REG = 2'b00,
  FU_SRC_MEM = 2'b01,
  FU_SRC_WB  = 2'b10
} fu_src_e;

typedef enum logic [1:0] {
  ALU_SRC_IMM,
  ALU_SRC_RS1,
  ALU_SRC_RS2
} alu_src_e;

typedef enum logic [2:0] {
  UNDEF,
  BYTE_S,
  BYTE_U,
  HALF_S,
  HALF_U,
  WORD
} data_size_e;