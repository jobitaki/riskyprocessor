package constants;
  parameter int ADDR_WIDTH = 9;
  parameter int SIM_MEM_SIZE = 16'hFFFF;

  typedef enum logic [31:0] {
    // I-type instructions
    I_LB        = 32'b????_????_????_????_?000_????_?000_0011,
    I_LH        = 32'b????_????_????_????_?001_????_?000_0011,
    I_LW        = 32'b????_????_????_????_?010_????_?000_0011,
    I_LBU       = 32'b????_????_????_????_?100_????_?000_0011,
    I_LHU       = 32'b????_????_????_????_?101_????_?000_0011,
    I_ALL_LOADS = 32'b????_????_????_????_????_????_?000_0011,

    I_ADDI  = 32'b????_????_????_????_?000_????_?001_0011,
    I_SLTI  = 32'b????_????_????_????_?010_????_?001_0011,
    I_SLTIU = 32'b????_????_????_????_?011_????_?001_0011,
    I_XORI  = 32'b????_????_????_????_?100_????_?001_0011,
    I_ORI   = 32'b????_????_????_????_?110_????_?001_0011,
    I_ANDI  = 32'b????_????_????_????_?111_????_?001_0011,
    I_SLLI  = 32'b0000_000?_????_????_?001_????_?001_0011,
    I_SRLI  = 32'b0000_000?_????_????_?101_????_?001_0011,
    I_SRAI  = 32'b0100_000?_????_????_?101_????_?001_0011,

    I_JALR = 32'b????_????_????_????_?000_????_?110_0111,

    // R-type instructions
    R_ADD     = 32'b0000_000?_????_????_?000_????_?011_0011,
    R_SUB     = 32'b0100_000?_????_????_?000_????_?011_0011,
    R_SLL     = 32'b0000_000?_????_????_?001_????_?011_0011,
    R_SLT     = 32'b0000_000?_????_????_?010_????_?011_0011,
    R_SLTU    = 32'b0000_000?_????_????_?011_????_?011_0011,
    R_XOR     = 32'b0000_000?_????_????_?100_????_?011_0011,
    R_SRL     = 32'b0000_000?_????_????_?101_????_?011_0011,
    R_SRA     = 32'b0100_000?_????_????_?101_????_?011_0011,
    R_OR      = 32'b0000_000?_????_????_?110_????_?011_0011,
    R_AND     = 32'b0000_000?_????_????_?111_????_?011_0011,
    R_ALL     = 32'b????_????_????_????_????_????_?011_0011,

    // S-type instructions
    S_SB  = 32'b????_????_????_????_?000_????_?010_0011, 
    S_SH  = 32'b????_????_????_????_?001_????_?010_0011, 
    S_SW  = 32'b????_????_????_????_?010_????_?010_0011,
    S_ALL = 32'b????_????_????_????_????_????_?010_0011,

    // B-type instructions
    B_BEQ  = 32'b????_????_????_????_?000_????_?110_0011,
    B_BNE  = 32'b????_????_????_????_?001_????_?110_0011,
    B_BLT  = 32'b????_????_????_????_?100_????_?110_0011,
    B_BGE  = 32'b????_????_????_????_?101_????_?110_0011,
    B_BLTU = 32'b????_????_????_????_?110_????_?110_0011,
    B_BGEU = 32'b????_????_????_????_?111_????_?110_0011,

    // J-type instructions
    J_JAL = 32'b????_????_????_????_????_????_?110_1111
    
  } opcode_e;

  typedef enum logic [3:0] {
    ALU_ADD   = 4'b0000,
    ALU_SUB   = 4'b0001,
    ALU_SLL   = 4'b0010,
    ALU_SLT   = 4'b0011,
    ALU_SLTU  = 4'b0100,
    ALU_XOR   = 4'b0101,
    ALU_SRL   = 4'b0110,
    ALU_SRA   = 4'b0111,
    ALU_OR    = 4'b1000,
    ALU_AND   = 4'b1001,
    ALU_NE    = 4'b1010,
    ALU_EQ    = 4'b1011,
    ALU_PASS  = 4'b1100,
    ALU_UNDEF = 4'b1111
  } alu_op_e;

  typedef enum logic [1:0] {
    FU_SRC_REG = 2'b00,
    FU_SRC_MEM = 2'b01,
    FU_SRC_WB  = 2'b10
  } fu_src_e;

  typedef enum logic [1:0] {
    ALU_SRC_IMM,
    ALU_SRC_RS1,
    ALU_SRC_RS2,
    ALU_SRC_PC
  } alu_src_e;

  typedef enum logic [2:0] {
    UNDEF,
    BYTE_S,
    BYTE_U,
    HALF_S,
    HALF_U,
    WORD
  } data_size_e;
endpackage